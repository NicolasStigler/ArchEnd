module condlogic (
  clk,
  reset,
  Cond,
  ALUFlags,
  FlagW,
  PCS,
  NextPC,
  RegW,
  MemW,
  PCWrite,
  RegWrite,
  MemWrite
);
  input wire clk;
  input wire reset;
  input wire [3:0] Cond;
  input wire [3:0] ALUFlags;
  input wire [1:0] FlagW;
  input wire PCS;
  input wire NextPC;
  input wire RegW;
  input wire MemW;
  output wire PCWrite;
  output wire RegWrite;
  output wire MemWrite;
  wire [1:0] FlagWrite;
  wire [3:0] Flags;
  wire CondEx;

  // Delay writing flags until ALUWB state
  flopr #(2) flagwritereg(
    clk,
    reset,
    FlagW & {2 {CondEx}},
    FlagWrite
  );

  // ADD CODE HERE

endmodule
